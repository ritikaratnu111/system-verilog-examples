// --------------------------------------------
// Design Name	:	parallel_fir
// File Name	:	types_and_constants.sv
// Function 	:	Package File for data types and constants
// Author	:	Ritika Ratnu
// ----------------------------------------------

package pkg;

	parameter SAMPLE_WIDTH	=	10;
	parameter FILTER_TAPS	=	13; 
endpackage: pkg

